    `timescale 1ns / 1ps

      module Infrarrojo(
      input [4:0] input_infra,
      output [4:0] output_infra
    );

     assign output_infra = input_infra;

    endmodule
